
// Verilog stimulus file.
// Please do not create a module in this file.


// Default verilog stimulus. 

initial
begin 

   cdsNet1 = 1'b0;
   cdsNet0 = 1'b0;
   io_VDD = 1'bz;
   io_VSS = 1'bz;
end 
