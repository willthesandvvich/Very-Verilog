// Global nets module 

`celldefine
module cds_globals;


supply0 gnd_;


endmodule
`endcelldefine
