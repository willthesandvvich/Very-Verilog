/home/seas/ugrad/tle14/ece468/ota_svrun1/ihnl/cds0/netlist